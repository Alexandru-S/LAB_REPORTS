-----------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;



entity mux_d is
end mux_d;

architecture Behavioral of mux_d is

begin


end Behavioral;

